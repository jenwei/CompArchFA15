module testFSM;

endmodule
