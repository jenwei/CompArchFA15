module ifu
(
output[31:0] 	instr,
input[25:0]	targetInstr,
input[15:0]	imm16,
input		branch,
input		jump
);
// controls/updates program counter
endmodule
