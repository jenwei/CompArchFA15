module testLUT;

endmodule
