module instrdec
(

);
// takes 32-bit instruction and outputs control signals
endmodule
