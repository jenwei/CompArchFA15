module cpu
(
);
// puts everything together 
// pulls instruction from register
// decodes instruction
// does things
ifu ifyou();
instrdecode ideeco();
fsm();



endmodule
