module testIFU;

endmodule
