module testSIGNEXTEND;

endmodule
