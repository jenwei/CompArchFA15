module cpu
(
input[31:0] instruction
);
// puts everything together =)
endmodule