module testDATAMEM;

endmodule
