module testMUX;

endmodule
