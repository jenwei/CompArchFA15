module instrdec
(
output jump,
output branch,

);
// takes 32-bit instruction and outputs control signals
endmodule
