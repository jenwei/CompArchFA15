module fsm
(

);
//Tracks state and controls enables
endmodule
