module testINSTRDEC;

endmodule
