module testCPU;

endmodule
