// Midpoint Check In
// -----------------

module midpoint(clk, sw, btn, led);
    input clk,
    input  [1:0] sw,
    input btn,
    output [3:0] led

endmodule
