module datamem
(
output[31:0]	dOut,
input[31:0] 	dIn,
input[31:0]	Addr,
input		memEnable
);
// Stores and retrieves program data
endmodule
