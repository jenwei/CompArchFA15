module regfile
(
output[31:0]	dA,
output[31:0]	dB,
input[31:0]	aA,
input[31:0]	aB,
input[31:0]	aW,
input[31:0]	dW,
input		wrEn
);
// tracks local data
endmodule