module testREGFILE;

endmodule
